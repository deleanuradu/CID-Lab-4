module top (input reg [1:0] in0,
				input reg [1:0] in1,		
				input reg sel,		
				output [3:0] out0,
		      output out1)

 out0 = 



				
						
endmodule						